library verilog;
use verilog.vl_types.all;
entity Sdram_Control_4Port is
    generic(
        INIT_PER        : integer := 24000;
        REF_PER         : integer := 1024;
        SC_CL           : integer := 3;
        SC_RCD          : integer := 3;
        SC_RRD          : integer := 7;
        SC_PM           : integer := 1;
        SC_BL           : integer := 1;
        SDR_BL          : vl_notype;
        SDR_BT          : vl_logic := Hi0;
        SDR_CL          : vl_notype
    );
    port(
        REF_CLK         : in     vl_logic;
        RESET_N         : in     vl_logic;
        CLK             : in     vl_logic;
        WR1_DATA        : in     vl_logic_vector(15 downto 0);
        WR1             : in     vl_logic;
        WR1_ADDR        : in     vl_logic_vector(22 downto 0);
        WR1_MAX_ADDR    : in     vl_logic_vector(22 downto 0);
        WR1_LENGTH      : in     vl_logic_vector(8 downto 0);
        WR1_LOAD        : in     vl_logic;
        WR1_CLK         : in     vl_logic;
        WR2_DATA        : in     vl_logic_vector(15 downto 0);
        WR2             : in     vl_logic;
        WR2_ADDR        : in     vl_logic_vector(22 downto 0);
        WR2_MAX_ADDR    : in     vl_logic_vector(22 downto 0);
        WR2_LENGTH      : in     vl_logic_vector(8 downto 0);
        WR2_LOAD        : in     vl_logic;
        WR2_CLK         : in     vl_logic;
        RD1_DATA        : out    vl_logic_vector(15 downto 0);
        RD1             : in     vl_logic;
        RD1_ADDR        : in     vl_logic_vector(22 downto 0);
        RD1_MAX_ADDR    : in     vl_logic_vector(22 downto 0);
        RD1_LENGTH      : in     vl_logic_vector(8 downto 0);
        RD1_LOAD        : in     vl_logic;
        RD1_CLK         : in     vl_logic;
        RD2_DATA        : out    vl_logic_vector(15 downto 0);
        RD2             : in     vl_logic;
        RD2_ADDR        : in     vl_logic_vector(22 downto 0);
        RD2_MAX_ADDR    : in     vl_logic_vector(22 downto 0);
        RD2_LENGTH      : in     vl_logic_vector(8 downto 0);
        RD2_LOAD        : in     vl_logic;
        RD2_CLK         : in     vl_logic;
        SA              : out    vl_logic_vector(11 downto 0);
        BA              : out    vl_logic_vector(1 downto 0);
        CS_N            : out    vl_logic_vector(1 downto 0);
        CKE             : out    vl_logic;
        RAS_N           : out    vl_logic;
        CAS_N           : out    vl_logic;
        WE_N            : out    vl_logic;
        DQ              : inout  vl_logic_vector(15 downto 0);
        DQM             : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of INIT_PER : constant is 1;
    attribute mti_svvh_generic_type of REF_PER : constant is 1;
    attribute mti_svvh_generic_type of SC_CL : constant is 1;
    attribute mti_svvh_generic_type of SC_RCD : constant is 1;
    attribute mti_svvh_generic_type of SC_RRD : constant is 1;
    attribute mti_svvh_generic_type of SC_PM : constant is 1;
    attribute mti_svvh_generic_type of SC_BL : constant is 1;
    attribute mti_svvh_generic_type of SDR_BL : constant is 3;
    attribute mti_svvh_generic_type of SDR_BT : constant is 1;
    attribute mti_svvh_generic_type of SDR_CL : constant is 3;
end Sdram_Control_4Port;
